		library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.filterpack.ALL;

entity FiltCte is
	port(
		ctes: out cte_t(N-1 downto 0)
		);
end FiltCte;

architecture arch of FiltCte is

begin

--Hamming 26 coeficientes precision 18 bits (1E-5)
--	ctes(0) <= "000000000011110110";
--	ctes(1) <= "000000000000011011";
--	ctes(2) <= "111111111000110001";
--	ctes(3) <= "111111110100000010";
--	ctes(4) <= "000000000001110001";
--	ctes(5) <= "000000011111111011";
--	ctes(6) <= "000000100110111100";
--	ctes(7) <= "111111101110101100";
--	ctes(8) <= "111110011000011101";
--	ctes(9) <= "111110011011010100";
--	ctes(10) <= "000001011010111100";
--	ctes(11) <= "000110100010110110";
--	ctes(12) <= "001010100110000101";
--	ctes(13) <= "001010100110000101";
--	ctes(14) <= "000110100010110110";
--	ctes(15) <= "000001011010111100";
--	ctes(16) <= "111110011011010100";
--	ctes(17) <= "111110011000011101";
--	ctes(18) <= "111111101110101100";
--	ctes(19) <= "000000100110111100";
--	ctes(20) <= "000000011111111011";
--	ctes(21) <= "000000000001110001";
--	ctes(22) <= "111111110100000010";
--	ctes(23) <= "111111111000110001";
--	ctes(24) <= "000000000000011011";
--	ctes(25) <= "000000000011110110";
	
--Hamming 26 coeficientes precision 21 bits (1E-6)
	ctes(0) <= "000000000011110110100";
	ctes(1) <= "000000000000011010111";
	ctes(2) <= "111111111000110000101";
	ctes(3) <= "111111110100000010011";
	ctes(4) <= "000000000001110000111";
	ctes(5) <= "000000011111111010110";
	ctes(6) <= "000000100110111100001";
	ctes(7) <= "111111101110101100010";
	ctes(8) <= "111110011000011100101";
	ctes(9) <= "111110011011010011111";
	ctes(10) <= "000001011010111011101";
	ctes(11) <= "000110100010110110001";
	ctes(12) <= "001010100110000101011";
	ctes(13) <= "001010100110000101011";
	ctes(14) <= "000110100010110110001";
	ctes(15) <= "000001011010111011101";
	ctes(16) <= "111110011011010011111";
	ctes(17) <= "111110011000011100101";
	ctes(18) <= "111111101110101100010";
	ctes(19) <= "000000100110111100001";
	ctes(20) <= "000000011111111010110";
	ctes(21) <= "000000000001110000111";
	ctes(22) <= "111111110100000010011";
	ctes(23) <= "111111111000110000101";
	ctes(24) <= "000000000000011010111";
	ctes(25) <= "000000000011110110100";
end arch;